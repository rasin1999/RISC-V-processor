module lsu(	input  [2:0] funct3,	output reg LoadType, StoreType);	always @(*)		case(funct3)			3'b000: {LoadType, StoreType} = 2'b01;			3'b010: {LoadType, StoreType} = 2'b00;			3'b100: {LoadType, StoreType} = 2'b1x;			default: {LoadType, StoreType} = 2'bxx;		endcaseendmodule